library ieee;
use ieee.std_logic_1164.all;

entity somadorHierarquico is
	port(A, B: in		std_logic_vector(n-1 downto 0)
			cin: in		std_logic;
			S: out		std_logic_vector(n-1 downto 0)
			
	)
end somadorHierarquico;